<svg xmlns="http://www.w3.org/2000/svg" width="180" height="36" viewBox="0 0 600 120">
  <defs>
    <linearGradient id="g" x1="0" y1="0" x2="1" y2="1">
      <stop offset="0" stop-color="#6ea8fe"/>
      <stop offset="1" stop-color="#88f0b2"/>
    </linearGradient>
  </defs>
  <rect width="600" height="120" fill="none"/>
  <text x="10" y="80" font-family="Montserrat,Segoe UI,Arial" font-size="72" font-weight="800" fill="url(#g)">AOMI</text>
  <text x="330" y="80" font-family="Montserrat,Segoe UI,Arial" font-size="48" font-weight="600" fill="#e8edf7" opacity=".9">Protocol</text>
</svg>
